/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  decoder.v                                          //
//                                                                     //
//  Description :  instruction decode (ID) stage of the pipeline;      // 
//                 decode the instruction fetch register operands, and // 
//                 compute immediate operand (if applicable)           // 
//                                                                     //
/////////////////////////////////////////////////////////////////////////


`timescale 1ns/100ps


  // Decode an instruction: given instruction bits IR produce the
  // appropriate datapath control signals.
  //
  // This is a *combinational* module (basically a PLA).
  //
module decoder(

	//input [31:0] inst,
	//input valid_inst_in,  // ignore inst when low, outputs will
	                      // reflect noop (except valid_inst)
	//see sys_defs.svh for definition
	input INST inst, 
	
	output ALU_OPA_SELECT opa_select,
	output ALU_OPB_SELECT opb_select,
	output DEST_REG_SEL   dest_reg, // mux selects
	output ALU_FUNC       alu_func,
	output FU_TYPE		  fu_type,
	output logic          is_jalr,
	output logic          rd_mem, wr_mem, cond_branch, uncond_branch,
	output MEM_SIZE       mem_size,
	output logic          load_signed,
	output logic          csr_op,    // used for CSR operations, we only used this as 
	                        //a cheap way to get the return code out
	output logic          halt,      // non-zero on a halt
	output logic          illegal,    // non-zero on an illegal instruction
	output logic          valid_inst  // for counting valid instructions executed
	                        // and for making the fetch stage die on halts/
	                        // keeping track of when to allow the next
	                        // instruction out of fetch
	                        // 0 for HALT and illegal instructions (die on halt)

); 
	assign valid_inst    =  ~illegal;
	always_comb begin
		// default control values:
		// - valid instructions must override these defaults as necessary.
		//	 opa_select, opb_select, and alu_func should be set explicitly.
		// - invalid instructions should clear valid_inst.
		// - These defaults are equivalent to a noop
		// * see sys_defs.vh for the constants used here
		opa_select = OPA_IS_RS1;
		opb_select = OPB_IS_RS2;
		alu_func = ALU_ADD;
		dest_reg = DEST_NONE;
		csr_op = `FALSE;
		rd_mem = `FALSE;
		wr_mem = `FALSE;
		cond_branch = `FALSE;
		uncond_branch = `FALSE;
		halt = `FALSE;
		illegal = `FALSE;
		fu_type = ALU;
		is_jalr = `FALSE;
		mem_size = WORD;
		load_signed = `FALSE;
		casez (inst) 
			`RV32_LUI: begin
				dest_reg   = DEST_RD;
				opa_select = OPA_IS_ZERO;
				opb_select = OPB_IS_U_IMM;
			end
			`RV32_AUIPC: begin
				dest_reg   = DEST_RD;
				opa_select = OPA_IS_PC;
				opb_select = OPB_IS_U_IMM;
			end
			`RV32_JAL: begin
				dest_reg      = DEST_RD;
				opa_select    = OPA_IS_PC;
				opb_select    = OPB_IS_J_IMM;
				uncond_branch = `TRUE;
				fu_type = BRANCH;
			end
			`RV32_JALR: begin
				dest_reg      = DEST_RD;
				opa_select    = OPA_IS_RS1;
				opb_select    = OPB_IS_I_IMM;
				uncond_branch = `TRUE;
				is_jalr       = `TRUE;
				fu_type = BRANCH;
			end
			`RV32_BEQ, `RV32_BNE, `RV32_BLT, `RV32_BGE,
			`RV32_BLTU, `RV32_BGEU: begin
				opa_select  = OPA_IS_PC;
				opb_select  = OPB_IS_B_IMM;
				cond_branch = `TRUE;
				fu_type = BRANCH;
			end
			`RV32_LB, `RV32_LH, `RV32_LW,
			`RV32_LBU, `RV32_LHU: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				rd_mem     = `TRUE;
				fu_type    = LOAD;
				mem_size   =  MEM_SIZE'(inst.r.funct3[1:0]);
				load_signed =	~inst.r.funct3[2];
			end
			`RV32_SB, `RV32_SH, `RV32_SW: begin
				opb_select = OPB_IS_S_IMM;
				wr_mem     = `TRUE;
				fu_type    = STORE;
				mem_size   =  MEM_SIZE'(inst.r.funct3[1:0]);
			end
			`RV32_ADDI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
			end
			`RV32_SLTI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_SLT;
			end
			`RV32_SLTIU: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_SLTU;
			end
			`RV32_ANDI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_AND;
			end
			`RV32_ORI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_OR;
			end
			`RV32_XORI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_XOR;
			end
			`RV32_SLLI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_SLL;
			end
			`RV32_SRLI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_SRL;
			end
			`RV32_SRAI: begin
				dest_reg   = DEST_RD;
				opb_select = OPB_IS_I_IMM;
				alu_func   = ALU_SRA;
			end
			`RV32_ADD: begin
				dest_reg   = DEST_RD;
			end
			`RV32_SUB: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_SUB;
			end
			`RV32_SLT: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_SLT;
			end
			`RV32_SLTU: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_SLTU;
			end
			`RV32_AND: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_AND;
			end
			`RV32_OR: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_OR;
			end
			`RV32_XOR: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_XOR;
			end
			`RV32_SLL: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_SLL;
			end
			`RV32_SRL: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_SRL;
			end
			`RV32_SRA: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_SRA;
			end
			`RV32_MUL: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_MUL;
				fu_type    = MUL;
			end
			`RV32_MULH: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_MULH;
				fu_type    = MUL;
			end
			`RV32_MULHSU: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_MULHSU;
				fu_type    = MUL;
			end
			`RV32_MULHU: begin
				dest_reg   = DEST_RD;
				alu_func   = ALU_MULHU;
				fu_type    = MUL;
			end
			`RV32_CSRRW, `RV32_CSRRS, `RV32_CSRRC: begin
				csr_op = `TRUE;
			end
			`WFI: begin
				halt = `TRUE;
			end
			default: illegal = `TRUE;
	endcase // casez (inst) 
	end // always
endmodule // decoder
 