//////////////////////////////////////////////////////////////////////////
//                                                                      //
//   Modulename :  rob.v                                                //                                                                     //
//  Description :  reorder buffer                                       //
//                                                                      // 
//////////////////////////////////////////////////////////////////////////


`define DEBUG
`ifndef __ROB_V__
`define __ROB_V__

`timescale 1ns/100ps

module rob(
    input                       clock,
    input                       reset,
    input [`XLEN-1:0]           PC,
    // dispatch
    input                       dispatch_enable,         // not only depend on rob_full, (e.g. invalid instr)
    input [4:0]                 dest_areg_idx,
    input [`PRF_LEN-1:0]        prf_free_preg_idx,
    input                       cond_branch,
    input                       uncond_branch,
    input                       local_pred_direction,
    input                       global_pred_direction,
    // cdb broadcast
    input                       cdb_broadcast_valid,     // make executed_rob_idx valid
    input [`ROB_LEN-1:0]        executed_rob_idx,                      
    input                       cdb_br_prediction,
    input                       cdb_br_target_PC,
    input                       cdb_mis_pred,

    //Outputs
    output logic [4:0]          rob_commit_dest_areg_idx,
    output logic [`PRF_LEN-1:0] rob_commit_dest_preg_idx,
    output logic [`ROB_LEN-1:0] rob_tail,
    output logic                rob_full,
    output logic                commit_valid,           // tell RRAT rob_commit_dest_(p|a)reg_idx is valid
    output logic [`XLEN-1:0]    result_PC,
    output logic                result_cond_branch,
    output logic                result_uncond_branch,
    output logic [`XLEN-1:0]    result_target_PC,
    output logic                result_local_pred_direction,
    output logic                result_global_pred_direction,
    output logic                result_branch_direction,
    output logic                mis_pred_is_head
);

    logic [`ROB_LEN-1:0]          rob_head;
    logic                         rob_empty;
    ROB_PACKET [`ROB_SIZE-1:0]    rob_packets;
     
    logic [`ROB_LEN:0]            rob_counter;

    assign commit_valid                 = (rob_packets[rob_head].executed) && (~rob_empty);
    assign rob_commit_dest_areg_idx     = rob_packets[rob_head].dest_areg_idx;
    assign rob_commit_dest_preg_idx     = rob_packets[rob_head].dest_preg_idx;
    assign rob_full                     = (rob_head == rob_tail) & (rob_counter != 0);
    assign result_PC                    = rob_packets[rob_head].PC;
    assign result_cond_branch           = rob_packets[rob_head].cond_branch;
    assign result_uncond_branch         = rob_packets[rob_head].uncond_branch;
    assign result_target_PC             = rob_packets[rob_head].target_PC;
    assign result_local_pred_direction  = rob_packets[rob_head].local_pred_direction;
    assign result_global_pred_direction = rob_packets[rob_head].global_pred_direction;
    assign result_branch_direction      = rob_packets[rob_head].branch_direction;
    assign mis_pred_is_head             = rob_packets[rob_head].rob_mis_pred && commit_valid;
    assign rob_empty                    = (rob_counter == 0);

    always_ff @(posedge clock) begin
        if (reset) begin
            rob_head    <= `SD `ROB_LEN'b0;
            rob_tail    <= `SD `ROB_LEN'b0; 
            rob_counter <= `SD `ROB_LEN'h0;
        end
        else if (mis_pred_is_head) begin
            rob_head    <= `SD rob_tail;
            rob_counter <= `SD `ROB_LEN'h0;
        end
        else begin 
            if (dispatch_enable) begin
                // dispatch
                rob_packets[rob_tail].PC                    <= `SD PC;
                rob_packets[rob_tail].executed              <= `SD 1'b0;
                rob_packets[rob_tail].dest_preg_idx         <= `SD prf_free_preg_idx;
                rob_packets[rob_tail].dest_areg_idx         <= `SD dest_areg_idx;
                rob_packets[rob_tail].rob_mis_pred          <= `SD 1'b0; 
                rob_packets[rob_tail].cond_branch           <= `SD cond_branch;
                rob_packets[rob_tail].uncond_branch         <= `SD uncond_branch;
                rob_packets[rob_tail].target_PC             <= `SD `XLEN'hfacebeec 
                rob_packets[rob_tail].local_pred_direction  <= `SD local_pred_direction;
                rob_packets[rob_tail].global_pred_direction <= `SD global_pred_direction;
                rob_packets[rob_tail].branch_direction      <= `SD 1'b0;
                rob_packets[rob_tail].branch_mis_pred       <= `SD cdb_mis_pred;
                rob_tail                                    <= `SD (rob_tail == `ROB_SIZE-1)? 0: rob_tail + 1;
            end  
            if(commit_valid) begin
                rob_head                            <= `SD (rob_head == `ROB_SIZE-1)? 0: rob_head + 1;
            end 
            if (cdb_broadcast_valid) begin
                //execute
                rob_packets[executed_rob_idx].executed         <= `SD 1'b1;
                rob_packets[executed_rob_idx].branch_direction <= `SD cdb_br_prediction;
                rob_packets[executed_rob_idx].target_PC        <= `Sd cdb_br_target_PC;
                rob_packets[executed_rob_idx].branch_mis_pred  <= `SD cdb_mis_pred;
            end
            rob_counter <= `SD (dispatch_enable && ~commit_valid) ? rob_counter+1 :
                               (~dispatch_enable && commit_valid) ? rob_counter-1 : rob_counter;

        end  
    end

endmodule
`endif // `__ROB_V__